module vlas

#flag linux -O2 -I/usr/local/include -I/usr/lib
#flag linux -L/usr/local/lib -L/usr/lib
#flag windows -O2
#flag windows -lgfortran
#flag darwin -I/usr/local/opt/lapacke/include
#flag darwin -L/usr/local/opt/lapacke/lib
#flag -I@VMODROOT
#flag -llapacke
