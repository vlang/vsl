module vsl

