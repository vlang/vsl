module fft

#flag linux -I/usr/local/include -I@VMODROOT
#flag linux -L/usr/lib -L/usr/local/lib
#flag darwin -I/usr/local/include -I@VMODROOT
#flag freebsd -I/usr/local/include -I@VMODROOT
#flag freebsd -L/usr/local/lib
#flag openbsd -I/usr/local/include -I@VMODROOT

#flag -lm
