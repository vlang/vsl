module native

#flag -I@VMODROOT

#include <vcl.h>
