module vcl

#flag linux -I@VMODROOT
#flag termux -I@VMODROOT
//#flag android -I@VMODROOT TODO try it
#flag windows -I@VMODROOT
#flag darwin -I@VMODROOT

#include <vcl.h>
