// Copyright (c) 2019 Ulises Jeremias Cornejo Fandos. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module specfunc

const (
        g                = 9.65657815377331589457187
        exp_g_o_sqrt_2pi = 6.23316569877722552586386e+3
        log_sqrt_2pi     = 9.18938533204672741780329736e-1


        gamma_a = [
                1.14400529453851095667309e+4,
                -3.23988020152318335053598e+4,
                3.50514523505571666566083e+4,
                -1.81641309541260702610647e+4,
                4.63232990536666818409138e+3,
                -5.36976777703356780555748e+2,
                2.28754473395181007645155e+1,
                -2.17925748738865115560082e-1,
                1.08314836272589368860689e-4
        ]


        /* Bernoulli numbers B(2),B(4),B(6),...,B(20).  Only B(2),...,B(6)
        * currently used.
        */

        B = [
                1.0 / f64(6 * 2 * 1),
                -1.0 / f64(30 * 4 * 3),
                1.0 / f64(42 * 6 * 5),
                -1.0 / f64(30 * 8 * 7),
                5.0 / f64(66 * 10 * 9),
                -691.0 / f64(2730 * 12 * 11),
                7.0 / f64(6 * 14 * 13),
                -3617.0 / f64(510 * 16 * 15),
                43867.0 / f64(796 * 18 * 17),
                -174611.0 / f64(330 * 20 * 19)
        ]
)
