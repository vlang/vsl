module blas
