module vcldl

import dl

pub const (
	default_paths = [
		'OpenCL${dl.dl_ext}',
	]
)
