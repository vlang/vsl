module vlas

import runtime
import sync
import vsl.blas.vlas.internal.float64
import vsl.util

