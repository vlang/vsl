module vsl
