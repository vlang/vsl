module dl

import dl

pub const (
	default_paths = [
		'OpenCL${dl.dl_ext}',
	]
)
