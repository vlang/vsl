// Copyright (c) 2019 Ulises Jeremias Cornejo Fandos. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module specfunc

const (
        eul = 0.57721566490153286061

        digamma_a = [
        f64(8.33333333333333333333e-2),
        -2.10927960927960927961e-2,
        7.57575757575757575758e-3,
        -4.16666666666666666667e-3,
        3.96825396825396825397e-3,
        -8.33333333333333333333e-3,
        8.33333333333333333333e-2
        ]
)
