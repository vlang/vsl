// Copyright (c) 2019-2020 Ulises Jeremias Cornejo Fandos. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module fun

const (
        // for x in [inf, 8]=1/[0,0.125]
        p0r8 = [
            f64(0.00000000000000000000e+00),  // 0x0000000000000000
                -7.03124999999900357484e-02, // 0xBFB1FFFFFFFFFD32
                -8.08167041275349795626e+00, // 0xC02029D0B44FA779
                -2.57063105679704847262e+02, // 0xC07011027B19E863
                -2.48521641009428822144e+03, // 0xC0A36A6ECD4DCAFC
                -5.25304380490729545272e+03, // 0xC0B4850B36CC643D
        ]
        p0s8 = [
            f64(1.16534364619668181717e+02), // 0x405D223307A96751
                3.83374475364121826715e+03, // 0x40ADF37D50596938
                4.05978572648472545552e+04, // 0x40E3D2BB6EB6B05F
                1.16752972564375915681e+05, // 0x40FC810F8F9FA9BD
                4.76277284146730962675e+04, // 0x40E741774F2C49DC
        ]

        // for x in [8,4.5454]=1/[0.125,0.22001]
        p0r5 = [
            f64(-1.14125464691894502584e-11), // 0xBDA918B147E495CC
                -7.03124940873599280078e-02, // 0xBFB1FFFFE69AFBC6
                -4.15961064470587782438e+00, // 0xC010A370F90C6BBF
                -6.76747652265167261021e+01, // 0xC050EB2F5A7D1783
                -3.31231299649172967747e+02, // 0xC074B3B36742CC63
                -3.46433388365604912451e+02, // 0xC075A6EF28A38BD7
        ]
        p0s5 = [
            f64(6.07539382692300335975e+01), // 0x404E60810C98C5DE
                1.05125230595704579173e+03, // 0x40906D025C7E2864
                5.97897094333855784498e+03, // 0x40B75AF88FBE1D60
                9.62544514357774460223e+03, // 0x40C2CCB8FA76FA38
                2.40605815922939109441e+03, // 0x40A2CC1DC70BE864
        ]

        // for x in [4.547,2.8571]=1/[0.2199,0.35001]
        p0r3 = [
            f64(-2.54704601771951915620e-09), // 0xBE25E1036FE1AA86
                -7.03119616381481654654e-02, // 0xBFB1FFF6F7C0E24B
                -2.40903221549529611423e+00, // 0xC00345B2AEA48074
                -2.19659774734883086467e+01, // 0xC035F74A4CB94E14
                -5.80791704701737572236e+01, // 0xC04D0A22420A1A45
                -3.14479470594888503854e+01, // 0xC03F72ACA892D80F
        ]
        p0s3 = [
            f64(3.58560338055209726349e+01), // 0x4041ED9284077DD3
                3.61513983050303863820e+02, // 0x40769839464A7C0E
                1.19360783792111533330e+03, // 0x4092A66E6D1061D6
                1.12799679856907414432e+03, // 0x40919FFCB8C39B7E
                1.73580930813335754692e+02, // 0x4065B296FC379081
        ]

        // for x in [2.8570,2]=1/[0.3499,0.5]
        p0r2 = [
            f64(-8.87534333032526411254e-08), // 0xBE77D316E927026D
                -7.03030995483624743247e-02, // 0xBFB1FF62495E1E42
                -1.45073846780952986357e+00, // 0xBFF736398A24A843
                -7.63569613823527770791e+00, // 0xC01E8AF3EDAFA7F3
                -1.11931668860356747786e+01, // 0xC02662E6C5246303
                -3.23364579351335335033e+00, // 0xC009DE81AF8FE70F
        ]
        p0s2 = [
            f64(2.22202997532088808441e+01), // 0x40363865908B5959
                1.36206794218215208048e+02, // 0x4061069E0EE8878F
                2.70470278658083486789e+02, // 0x4070E78642EA079B
                1.53875394208320329881e+02, // 0x40633C033AB6FAFF
                1.46576176948256193810e+01, // 0x402D50B344391809
        ]

        // for x in [inf, 8]=1/[0,0.125]
        p1r8 = [
            f64(0.00000000000000000000e+00), // 0x0000000000000000
                1.17187499999988647970e-01, // 0x3FBDFFFFFFFFFCCE
                1.32394806593073575129e+01, // 0x402A7A9D357F7FCE
                4.12051854307378562225e+02, // 0x4079C0D4652EA590
                3.87474538913960532227e+03, // 0x40AE457DA3A532CC
                7.91447954031891731574e+03, // 0x40BEEA7AC32782DD
        ]
        p1s8 = [
            f64(1.14207370375678408436e+02), // 0x405C8D458E656CAC
                3.65093083420853463394e+03, // 0x40AC85DC964D274F
                3.69562060269033463555e+04, // 0x40E20B8697C5BB7F
                9.76027935934950801311e+04, // 0x40F7D42CB28F17BB
                3.08042720627888811578e+04, // 0x40DE1511697A0B2D
        ]

        // for x in [8,4.5454] = 1/[0.125,0.22001]
        p1r5 = [
            f64(1.31990519556243522749e-11), // 0x3DAD0667DAE1CA7D
                1.17187493190614097638e-01, // 0x3FBDFFFFE2C10043
                6.80275127868432871736e+00, // 0x401B36046E6315E3
                1.08308182990189109773e+02, // 0x405B13B9452602ED
                5.17636139533199752805e+02, // 0x40802D16D052D649
                5.28715201363337541807e+02, // 0x408085B8BB7E0CB7
        ]
        p1s5 = [
            f64(5.92805987221131331921e+01), // 0x404DA3EAA8AF633D
                9.91401418733614377743e+02, // 0x408EFB361B066701
                5.35326695291487976647e+03, // 0x40B4E9445706B6FB
                7.84469031749551231769e+03, // 0x40BEA4B0B8A5BB15
                1.50404688810361062679e+03, // 0x40978030036F5E51
        ]

        // for x in[4.5453,2.8571] = 1/[0.2199,0.35001]
        p1r3 = [
            f64(3.02503916137373618024e-09), // 0x3E29FC21A7AD9EDD
                1.17186865567253592491e-01, // 0x3FBDFFF55B21D17B
                3.93297750033315640650e+00, // 0x400F76BCE85EAD8A
                3.51194035591636932736e+01, // 0x40418F489DA6D129
                9.10550110750781271918e+01, // 0x4056C3854D2C1837
                4.85590685197364919645e+01, // 0x4048478F8EA83EE5
        ]
        p1s3 = [
            f64(3.47913095001251519989e+01), // 0x40416549A134069C
                3.36762458747825746741e+02, // 0x40750C3307F1A75F
                1.04687139975775130551e+03, // 0x40905B7C5037D523
                8.90811346398256432622e+02, // 0x408BD67DA32E31E9
                1.03787932439639277504e+02, // 0x4059F26D7C2EED53
        ]

        // for x in [2.8570,2] = 1/[0.3499,0.5]
        p1r2 = [
            f64(1.07710830106873743082e-07), // 0x3E7CE9D4F65544F4
                1.17176219462683348094e-01, // 0x3FBDFF42BE760D83
                2.36851496667608785174e+00, // 0x4002F2B7F98FAEC0
                1.22426109148261232917e+01, // 0x40287C377F71A964
                1.76939711271687727390e+01, // 0x4031B1A8177F8EE2
                5.07352312588818499250e+00, // 0x40144B49A574C1FE
        ]
        p1s2 = [
            f64(2.14364859363821409488e+01), // 0x40356FBD8AD5ECDC
                1.25290227168402751090e+02, // 0x405F529314F92CD5
                2.32276469057162813669e+02, // 0x406D08D8D5A2DBD9
                1.17679373287147100768e+02, // 0x405D6B7ADA1884A9
                8.36463893371618283368e+00, // 0x4020BAB1F44E5192
        ]

        // for x in [inf, 8]=1/[0,0.125]
        q0r8 = [
            f64(0.00000000000000000000e+00), // 0x0000000000000000
                7.32421874999935051953e-02, // 0x3FB2BFFFFFFFFE2C
                1.17682064682252693899e+01, // 0x402789525BB334D6
                5.57673380256401856059e+02, // 0x40816D6315301825
                8.85919720756468632317e+03, // 0x40C14D993E18F46D
                3.70146267776887834771e+04, // 0x40E212D40E901566
        ]
        q0s8 = [
            f64(1.63776026895689824414e+02),  // 0x406478D5365B39BC
                8.09834494656449805916e+03,  // 0x40BFA2584E6B0563
                1.42538291419120476348e+05,  // 0x4101665254D38C3F
                8.03309257119514397345e+05,  // 0x412883DA83A52B43
                8.40501579819060512818e+05,  // 0x4129A66B28DE0B3D
                -3.43899293537866615225e+05, // 0xC114FD6D2C9530C5
        ]

        // for x in [8,4.5454]=1/[0.125,0.22001]
        q0r5 = [
            f64(1.84085963594515531381e-11), // 0x3DB43D8F29CC8CD9
                7.32421766612684765896e-02, // 0x3FB2BFFFD172B04C
                5.83563508962056953777e+00, // 0x401757B0B9953DD3
                1.35111577286449829671e+02, // 0x4060E3920A8788E9
                1.02724376596164097464e+03, // 0x40900CF99DC8C481
                1.98997785864605384631e+03, // 0x409F17E953C6E3A6
        ]
        q0s5 = [
            f64(8.27766102236537761883e+01),  // 0x4054B1B3FB5E1543
                2.07781416421392987104e+03,  // 0x40A03BA0DA21C0CE
                1.88472887785718085070e+04,  // 0x40D267D27B591E6D
                5.67511122894947329769e+04,  // 0x40EBB5E397E02372
                3.59767538425114471465e+04,  // 0x40E191181F7A54A0
                -5.35434275601944773371e+03, // 0xC0B4EA57BEDBC609
        ]

        // for x in [4.547,2.8571]=1/[0.2199,0.35001]
        q0r3 = [
            f64(4.37741014089738620906e-09), // 0x3E32CD036ADECB82
                7.32411180042911447163e-02, // 0x3FB2BFEE0E8D0842
                3.34423137516170720929e+00, // 0x400AC0FC61149CF5
                4.26218440745412650017e+01, // 0x40454F98962DAEDD
                1.70808091340565596283e+02, // 0x406559DBE25EFD1F
                1.66733948696651168575e+02, // 0x4064D77C81FA21E0
        ]
        q0s3 = [
            f64(4.87588729724587182091e+01),  // 0x40486122BFE343A6
                7.09689221056606015736e+02,  // 0x40862D8386544EB3
                3.70414822620111362994e+03,  // 0x40ACF04BE44DFC63
                6.46042516752568917582e+03,  // 0x40B93C6CD7C76A28
                2.51633368920368957333e+03,  // 0x40A3A8AAD94FB1C0
                -1.49247451836156386662e+02, // 0xC062A7EB201CF40F
        ]

        // for x in [2.8570,2]=1/[0.3499,0.5]
        q0r2 = [
            f64(1.50444444886983272379e-07), // 0x3E84313B54F76BDB
                7.32234265963079278272e-02, // 0x3FB2BEC53E883E34
                1.99819174093815998816e+00, // 0x3FFFF897E727779C
                1.44956029347885735348e+01, // 0x402CFDBFAAF96FE5
                3.16662317504781540833e+01, // 0x403FAA8E29FBDC4A
                1.62527075710929267416e+01, // 0x403040B171814BB4
        ]
        q0s2 = [
            f64(3.03655848355219184498e+01),  // 0x403E5D96F7C07AED
                2.69348118608049844624e+02,  // 0x4070D591E4D14B40
                8.44783757595320139444e+02,  // 0x408A664522B3BF22
                8.82935845112488550512e+02,  // 0x408B977C9C5CC214
                2.12666388511798828631e+02,  // 0x406A95530E001365
                -5.31095493882666946917e+00, // 0xC0153E6AF8B32931
        ]

        // for x in [inf, 8] = 1/[0,0.125]
        q1r8 = [
            f64(0.00000000000000000000e+00),  // 0x0000000000000000
                -1.02539062499992714161e-01, // 0xBFBA3FFFFFFFFDF3
                -1.62717534544589987888e+01, // 0xC0304591A26779F7
                -7.59601722513950107896e+02, // 0xC087BCD053E4B576
                -1.18498066702429587167e+04, // 0xC0C724E740F87415
                -4.84385124285750353010e+04, // 0xC0E7A6D065D09C6A
        ]
        q1s8 = [
            f64(1.61395369700722909556e+02),  // 0x40642CA6DE5BCDE5
                7.82538599923348465381e+03,  // 0x40BE9162D0D88419
                1.33875336287249578163e+05,  // 0x4100579AB0B75E98
                7.19657723683240939863e+05,  // 0x4125F65372869C19
                6.66601232617776375264e+05,  // 0x412457D27719AD5C
                -2.94490264303834643215e+05, // 0xC111F9690EA5AA18
        ]

        // for x in [8,4.5454] = 1/[0.125,0.22001]
        q1r5 = [
            f64(-2.08979931141764104297e-11), // 0xBDB6FA431AA1A098
                -1.02539050241375426231e-01, // 0xBFBA3FFFCB597FEF
                -8.05644828123936029840e+00, // 0xC0201CE6CA03AD4B
                -1.83669607474888380239e+02, // 0xC066F56D6CA7B9B0
                -1.37319376065508163265e+03, // 0xC09574C66931734F
                -2.61244440453215656817e+03, // 0xC0A468E388FDA79D
        ]
        q1s5 = [
            f64(8.12765501384335777857e+01),  // 0x405451B2FF5A11B2
                1.99179873460485964642e+03,  // 0x409F1F31E77BF839
                1.74684851924908907677e+04,  // 0x40D10F1F0D64CE29
                4.98514270910352279316e+04,  // 0x40E8576DAABAD197
                2.79480751638918118260e+04,  // 0x40DB4B04CF7C364B
                -4.71918354795128470869e+03, // 0xC0B26F2EFCFFA004
        ]

        // for x in [4.5454,2.8571] = 1/[0.2199,0.35001] ???
        q1r3 = [
            f64(-5.07831226461766561369e-09), // 0xBE35CFA9D38FC84F
                -1.02537829820837089745e-01, // 0xBFBA3FEB51AEED54
                -4.61011581139473403113e+00, // 0xC01270C23302D9FF
                -5.78472216562783643212e+01, // 0xC04CEC71C25D16DA
                -2.28244540737631695038e+02, // 0xC06C87D34718D55F
                -2.19210128478909325622e+02, // 0xC06B66B95F5C1BF6
        ]
        q1s3 = [
            f64(4.76651550323729509273e+01),  // 0x4047D523CCD367E4
                6.73865112676699709482e+02,  // 0x40850EEBC031EE3E
                3.38015286679526343505e+03,  // 0x40AA684E448E7C9A
                5.54772909720722782367e+03,  // 0x40B5ABBAA61D54A6
                1.90311919338810798763e+03,  // 0x409DBC7A0DD4DF4B
                -1.35201191444307340817e+02, // 0xC060E670290A311F
        ]

        // for x in [2.8570,2] = 1/[0.3499,0.5]
        q1r2 = [
            f64(-1.78381727510958865572e-07), // 0xBE87F12644C626D2
                -1.02517042607985553460e-01, // 0xBFBA3E8E9148B010
                -2.75220568278187460720e+00, // 0xC006048469BB4EDA
                -1.96636162643703720221e+01, // 0xC033A9E2C168907F
                -4.23253133372830490089e+01, // 0xC04529A3DE104AAA
                -2.13719211703704061733e+01, // 0xC0355F3639CF6E52
        ]
        q1s2 = [
            f64(2.95333629060523854548e+01),  // 0x403D888A78AE64FF
                2.52981549982190529136e+02,  // 0x406F9F68DB821CBA
                7.57502834868645436472e+02,  // 0x4087AC05CE49A0F7
                7.39393205320467245656e+02,  // 0x40871B2548D4C029
                1.55949003336666123687e+02,  // 0x40637E5E3C3ED8D4
                -4.95949898822628210127e+00, // 0xC013D686E71BE86B
        ]
)
