// Copyright (c) 2019 Ulises Jeremias Cornejo Fandos. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.

module specfunc

const (
        log_sqrt_2pi = 9.18938533204672741780329736e-1

        B = [
        /* Bernoulli numbers B(2),B(4),B(6),...,B(20).  Only B(2),...,B(10) currently
        * used.
        */
    f64(1.0 / (6.0 * 2.0 * 1.0)),
       -1.0 / (30.0 * 4.0 * 3.0),
        1.0 / (42.0 * 6.0 * 5.0),
       -1.0 / (30.0 * 8.0 * 7.0),
        5.0 / (66.0 * 10.0 * 9.0),
       -691.0 / (2730.0 * 12.0 * 11.0),
        7.0 / (6.0 * 14.0 * 13.0),
       -3617.0 / (510.0 * 16.0 * 15.0),
        43867.0 / (796.0 * 18.0 * 17.0),
       -174611.0 / (330.0 * 20.0 * 19.0)
        ]


	log_factorials = [
    f64(0.000000000000000000000e+0),      /*   0! */
	0.000000000000000000000e+0,       /*   1! */
	6.931471805599453094172e-1,       /*   2! */
	1.791759469228055000812e+0,       /*   3! */
	3.178053830347945619647e+0,       /*   4! */
	4.787491742782045994248e+0,       /*   5! */
	6.579251212010100995060e+0,       /*   6! */
	8.525161361065414300166e+0,       /*   7! */
	1.060460290274525022842e+1,       /*   8! */
	1.280182748008146961121e+1,       /*   9! */
	1.510441257307551529523e+1,       /*  10! */
	1.750230784587388583929e+1,       /*  11! */
	1.998721449566188614952e+1,       /*  12! */
	2.255216385312342288557e+1,       /*  13! */
	2.519122118273868150009e+1,       /*  14! */
	2.789927138384089156609e+1,       /*  15! */
	3.067186010608067280376e+1,       /*  16! */
	3.350507345013688888401e+1,       /*  17! */
	3.639544520803305357622e+1,       /*  18! */
	3.933988418719949403622e+1,       /*  19! */
	4.233561646075348502966e+1,       /*  20! */
	4.538013889847690802616e+1,       /*  21! */
	4.847118135183522387964e+1,       /*  22! */
	5.160667556776437357045e+1,       /*  23! */
	5.478472939811231919009e+1,       /*  24! */
	5.800360522298051993929e+1,       /*  25! */
	6.126170176100200198477e+1,       /*  26! */
	6.455753862700633105895e+1,       /*  27! */
	6.788974313718153498289e+1,       /*  28! */
	7.125703896716800901007e+1,       /*  29! */
	7.465823634883016438549e+1,       /*  30! */
	7.809222355331531063142e+1,       /*  31! */
	8.155795945611503717850e+1,       /*  32! */
	8.505446701758151741396e+1,       /*  33! */
	8.858082754219767880363e+1,       /*  34! */
	9.213617560368709248333e+1,       /*  35! */
	9.571969454214320248496e+1,       /*  36! */
	9.933061245478742692933e+1,       /*  37! */
	1.029681986145138126988e+2,       /*  38! */
	1.066317602606434591262e+2,       /*  39! */
	1.103206397147573954291e+2,       /*  40! */
	1.140342117814617032329e+2,       /*  41! */
	1.177718813997450715388e+2,       /*  42! */
	1.215330815154386339623e+2,       /*  43! */
	1.253172711493568951252e+2,       /*  44! */
	1.291239336391272148826e+2,       /*  45! */
	1.329525750356163098828e+2,       /*  46! */
	1.368027226373263684696e+2,       /*  47! */
	1.406739236482342593987e+2,       /*  48! */
	1.445657439463448860089e+2,       /*  49! */
	1.484777669517730320675e+2,       /*  50! */
	1.524095925844973578392e+2,       /*  51! */
	1.563608363030787851941e+2,       /*  52! */
	1.603311282166309070282e+2,       /*  53! */
	1.643201122631951814118e+2,       /*  54! */
	1.683274454484276523305e+2,       /*  55! */
	1.723527971391628015638e+2,       /*  56! */
	1.763958484069973517152e+2,       /*  57! */
	1.804562914175437710518e+2,       /*  58! */
	1.845338288614494905025e+2,       /*  59! */
	1.886281734236715911873e+2,       /*  60! */
	1.927390472878449024360e+2,       /*  61! */
	1.968661816728899939914e+2,       /*  62! */
	2.010093163992815266793e+2,       /*  63! */
	2.051681994826411985358e+2,       /*  64! */
	2.093425867525368356464e+2,       /*  65! */
	2.135322414945632611913e+2,       /*  66! */
	2.177369341139542272510e+2,       /*  67! */
	2.219564418191303339501e+2,       /*  68! */
	2.261905483237275933323e+2,       /*  69! */
	2.304390435657769523214e+2,       /*  70! */
	2.347017234428182677427e+2,       /*  71! */
	2.389783895618343230538e+2,       /*  72! */
	2.432688490029827141829e+2,       /*  73! */
	2.475729140961868839366e+2,       /*  74! */
	2.518904022097231943772e+2,       /*  75! */
	2.562211355500095254561e+2,       /*  76! */
	2.605649409718632093053e+2,       /*  77! */
	2.649216497985528010421e+2,       /*  78! */
	2.692910976510198225363e+2,       /*  79! */
	2.736731242856937041486e+2,       /*  80! */
	2.780675734403661429141e+2,       /*  81! */
	2.824742926876303960274e+2,       /*  82! */
	2.868931332954269939509e+2,       /*  83! */
	2.913239500942703075662e+2,       /*  84! */
	2.957666013507606240211e+2,       /*  85! */
	3.002209486470141317540e+2,       /*  86! */
	3.046868567656687154726e+2,       /*  87! */
	3.091641935801469219449e+2,       /*  88! */
	3.136528299498790617832e+2,       /*  89! */
	3.181526396202093268500e+2,       /*  90! */
	3.226634991267261768912e+2,       /*  91! */
	3.271852877037752172008e+2,       /*  92! */
	3.317178871969284731381e+2,       /*  93! */
	3.362611819791984770344e+2,       /*  94! */
	3.408150588707990178690e+2,       /*  95! */
	3.453794070622668541074e+2,       /*  96! */
	3.499541180407702369296e+2,       /*  97! */
	3.545390855194408088492e+2,       /*  98! */
	3.591342053695753987760e+2,       /*  99! */
	3.637393755555634901441e+2,       /* 100! */
	3.683544960724047495950e+2,       /* 101! */
	3.729794688856890206760e+2,       /* 102! */
	3.776141978739186564468e+2,       /* 103! */
	3.822585887730600291111e+2,       /* 104! */
	3.869125491232175524822e+2,       /* 105! */
	3.915759882173296196258e+2,       /* 106! */
	3.962488170517915257991e+2,       /* 107! */
	4.009309482789157454921e+2,       /* 108! */
	4.056222961611448891925e+2,       /* 109! */
	4.103227765269373054205e+2,       /* 110! */
	4.150323067282496395563e+2,       /* 111! */
	4.197508055995447340991e+2,       /* 112! */
	4.244781934182570746677e+2,       /* 113! */
	4.292143918666515701285e+2,       /* 114! */
	4.339593239950148201939e+2,       /* 115! */
	4.387129141861211848399e+2,       /* 116! */
	4.434750881209189409588e+2,       /* 117! */
	4.482457727453846057188e+2,       /* 118! */
	4.530248962384961351041e+2,       /* 119! */
	4.578123879812781810984e+2,       /* 120! */
	4.626081785268749221865e+2,       /* 121! */
	4.674121995716081787447e+2,       /* 122! */
	4.722243839269805962399e+2,       /* 123! */
	4.770446654925856331047e+2,       /* 124! */
	4.818729792298879342285e+2,       /* 125! */
	4.867092611368394122258e+2,       /* 126! */
	4.915534482232980034989e+2,       /* 127! */
	4.964054784872176206648e+2,       /* 128! */
	5.012652908915792927797e+2,       /* 129! */
	5.061328253420348751997e+2,       /* 130! */
	5.110080226652360267439e+2,       /* 131! */
	5.158908245878223975982e+2,       /* 132! */
	5.207811737160441513633e+2,       /* 133! */
	5.256790135159950627324e+2,       /* 134! */
	5.305842882944334921812e+2,       /* 135! */
	5.354969431801695441897e+2,       /* 136! */
	5.404169241059976691050e+2,       /* 137! */
	5.453441777911548737966e+2,       /* 138! */
	5.502786517242855655538e+2,       /* 139! */
	5.552202941468948698523e+2,       /* 140! */
	5.601690540372730381305e+2,       /* 141! */
	5.651248810948742988613e+2,       /* 142! */
	5.700877257251342061414e+2,       /* 143! */
	5.750575390247102067619e+2,       /* 144! */
	5.800342727671307811636e+2,       /* 145! */
	5.850178793888391176022e+2,       /* 146! */
	5.900083119756178539038e+2,       /* 147! */
	5.950055242493819689670e+2,       /* 148! */
	6.000094705553274281080e+2,       /* 149! */
	6.050201058494236838580e+2,       /* 150! */
	6.100373856862386081868e+2,       /* 151! */
	6.150612662070848845750e+2,       /* 152! */
	6.200917041284773200381e+2,       /* 153! */
	6.251286567308909491967e+2,       /* 154! */
	6.301720818478101958172e+2,       /* 155! */
	6.352219378550597328635e+2,       /* 156! */
	6.402781836604080409209e+2,       /* 157! */
	6.453407786934350077245e+2,       /* 158! */
	6.504096828956552392500e+2,       /* 159! */
	6.554848567108890661717e+2,       /* 160! */
	6.605662610758735291676e+2,       /* 161! */
	6.656538574111059132426e+2,       /* 162! */
	6.707476076119126755767e+2,       /* 163! */
	6.758474740397368739994e+2,       /* 164! */
	6.809534195136374546094e+2,       /* 165! */
	6.860654073019939978423e+2,       /* 166! */
	6.911834011144107529496e+2,       /* 167! */
	6.963073650938140118743e+2,       /* 168! */
	7.014372638087370853465e+2,       /* 169! */
	7.065730622457873471107e+2,       /* 170! */
	7.117147258022900069535e+2,       /* 171! */
	]
)
