module plot

pub struct Font {
pub mut:
	color		string	= 'black'
	family		string	= 'monospace'
	size		f64		= 16.
	// WIP: new properties will be added eventually.
}
