module vcl


