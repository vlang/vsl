// Copyright (c) 2024. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module lapack

import math
import vsl.blas
import vsl.float.float64
import rand

// Test tolerance similar to gonum's LAPACK tests
const test_tolerance = 1e-12
const ortho_tolerance = 1e-15

// Test utilities and helpers

// nearly_equal_matrix checks if two matrices are nearly equal within tolerance
fn nearly_equal_matrix(a [][]f64, b [][]f64, tol f64) bool {
	dump('nearly_equal_matrix: a.len=${a.len}, b.len=${b.len}')
	if a.len != b.len {
		return false
	}
	for i in 0 .. a.len {
		dump('nearly_equal_matrix loop i=${i}: a[i].len=${a[i].len}, b[i].len=${b[i].len}')
		if a[i].len != b[i].len {
			return false
		}
		for j in 0 .. a[i].len {
			dump('nearly_equal_matrix: i=${i}, j=${j}, a[i].len=${a[i].len}')
			if !float64.tolerance(a[i][j], b[i][j], tol) {
				return false
			}
		}
	}
	return true
}

// matrix_norm computes various matrix norms
fn matrix_norm(a [][]f64, norm_type string) f64 {
	m := a.len
	if m == 0 {
		return 0.0
	}
	n := a[0].len
	if n == 0 {
		return 0.0
	}

	match norm_type {
		'fro' { // Frobenius norm
			mut sum := 0.0
			for i in 0 .. m {
				for j in 0 .. n {
					sum += a[i][j] * a[i][j]
				}
			}
			return math.sqrt(sum)
		}
		'1' { // 1-norm (maximum column sum)
			mut max_sum := 0.0
			for j in 0 .. n {
				mut col_sum := 0.0
				for i in 0 .. m {
					col_sum += math.abs(a[i][j])
				}
				if col_sum > max_sum {
					max_sum = col_sum
				}
			}
			return max_sum
		}
		'inf' { // infinity norm (maximum row sum)
			mut max_sum := 0.0
			for i in 0 .. m {
				mut row_sum := 0.0
				for j in 0 .. n {
					row_sum += math.abs(a[i][j])
				}
				if row_sum > max_sum {
					max_sum = row_sum
				}
			}
			return max_sum
		}
		else {
			return 0.0
		}
	}
}

// create_identity creates an n x n identity matrix
fn create_identity(n int) [][]f64 {
	mut id := [][]f64{len: n, init: []f64{len: n, init: 0.0}}
	for i in 0 .. n {
		id[i][i] = 1.0
	}
	return id
}

// create_random_matrix creates an m x n matrix with random values between -1 and 1
fn create_random_matrix(m int, n int, seed int) [][]f64 {
	rand.seed([u32(seed), u32(seed)])
	mut mat := [][]f64{len: m, init: []f64{len: n}}
	for i in 0 .. m {
		for j in 0 .. n {
			mat[i][j] = rand.f64_in_range(-1.0, 1.0) or { 0.0 }
		}
	}
	return mat
}

// create_spd_matrix creates a symmetric positive definite matrix for testing Cholesky
fn create_spd_matrix(n int, seed int) [][]f64 {
	// Create a random matrix and compute A'A to make it SPD
	a := create_random_matrix(n, n, seed)
	mut spd := [][]f64{len: n, init: []f64{len: n, init: 0.0}}

	// Compute A'A
	for i in 0 .. n {
		for j in 0 .. n {
			for k in 0 .. n {
				spd[i][j] += a[k][i] * a[k][j]
			}
		}
	}

	// Add some to diagonal for numerical stability
	for i in 0 .. n {
		spd[i][i] += 1.0
	}

	return spd
}

// matrix_multiply multiplies two matrices A and B
fn matrix_multiply(a [][]f64, b [][]f64) [][]f64 {
	m := a.len
	n := b[0].len
	k := a[0].len

	mut c := [][]f64{len: m, init: []f64{len: n, init: 0.0}}

	for i in 0 .. m {
		for j in 0 .. n {
			for l in 0 .. k {
				c[i][j] += a[i][l] * b[l][j]
			}
		}
	}
	return c
}

// matrix_transpose transposes a matrix
fn matrix_transpose(a [][]f64) [][]f64 {
	m := a.len
	n := a[0].len
	mut at := [][]f64{len: n, init: []f64{len: m}}

	for i in 0 .. m {
		for j in 0 .. n {
			at[j][i] = a[i][j]
		}
	}
	return at
}

// check_orthogonal verifies that a matrix has orthonormal columns/rows
fn check_orthogonal(q [][]f64, check_columns bool) bool {
	m := q.len
	n := q[0].len

	if check_columns {
		// Check Q'Q = I
		qt := matrix_transpose(q)
		qtq := matrix_multiply(qt, q)
		identity := create_identity(n)
		return nearly_equal_matrix(qtq, identity, ortho_tolerance)
	} else {
		// Check QQ' = I
		qqt := matrix_multiply(q, matrix_transpose(q))
		identity := create_identity(m)
		return nearly_equal_matrix(qqt, identity, ortho_tolerance)
	}
}

// ============================================================================
// GESV Tests - General Linear System Solver
// ============================================================================

fn test_gesv_basic() {
	// Test 1: Simple 2x2 system
	mut a := [[2.0, 1.0], [1.0, 1.0]]
	mut b := [[3.0, 5.0], [2.0, 3.0]] // Two RHS vectors

	original_a := a.clone()
	expected_x := [[1.0, 2.0], [1.0, 1.0]] // Known solution: Column 1: [1,1], Column 2: [2,1]

	gesv(mut a, mut b) or { assert false, 'gesv failed on simple 2x2 system' }

	// Check solution
	assert nearly_equal_matrix(b, expected_x, test_tolerance), 'gesv solution incorrect for 2x2 system'

	// Test 2: Verify by substitution: A * X = B (original)
	result := matrix_multiply(original_a, b)
	original_b := [[3.0, 5.0], [2.0, 3.0]]
	assert nearly_equal_matrix(result, original_b, test_tolerance), 'gesv: A*X != B'
}

fn test_gesv_square_systems() {
	// Test various sizes following gonum patterns
	sizes := [1, 3, 5, 10, 20]

	for n in sizes {
		// Create well-conditioned system
		mut a := create_identity(n)
		// Add some off-diagonal elements to make it non-trivial
		for i in 0 .. n - 1 {
			a[i][i + 1] = 0.5
			a[i + 1][i] = 0.3
		}

		// Create exact solution
		x_exact := create_random_matrix(n, 2, 42 + n) // 2 RHS vectors

		// Compute RHS: b = A * x_exact
		mut b := matrix_multiply(a, x_exact)

		// Solve the system
		mut a_copy := a.clone()
		gesv(mut a_copy, mut b) or { assert false, 'gesv failed for n=${n}' }

		// Check solution accuracy
		assert nearly_equal_matrix(b, x_exact, test_tolerance), 'gesv solution incorrect for n=${n}'

		// Verify residual: ||A*x - b_original|| should be small
		mut residual := matrix_multiply(a, b)
		b_original := matrix_multiply(a, x_exact)
		for i in 0 .. n {
			for j in 0 .. 2 {
				residual[i][j] -= b_original[i][j]
			}
		}
		residual_norm := matrix_norm(residual, 'fro')
		assert residual_norm < test_tolerance, 'gesv residual too large for n=${n}: ${residual_norm}'
	}
}

// ============================================================================
// GETRF/GETRI Tests - LU Factorization and Matrix Inversion
// ============================================================================

fn test_getrf_basic() {
	// Test 1: Simple 3x3 matrix
	mut a := [[2.0, 1.0, 1.0], [4.0, 3.0, 3.0], [8.0, 7.0, 9.0]]

	original_a := a.clone()

	ipiv := getrf(mut a) or {
		assert false, 'getrf failed on 3x3 matrix'
		return
	}

	// Check that pivot array has correct length and valid indices
	assert ipiv.len == 3, 'getrf: wrong pivot array length'
	for i, p in ipiv {
		assert p >= i && p < 3, 'getrf: invalid pivot index ${p} at position ${i}'
	}

	// Test 2: Verify LU factorization by reconstruction
	// Extract L and U from the result
	n := 3
	mut l := [][]f64{len: n, init: []f64{len: n, init: 0.0}}
	mut u := [][]f64{len: n, init: []f64{len: n, init: 0.0}}

	for i in 0 .. n {
		l[i][i] = 1.0 // L has unit diagonal
		for j in 0 .. i {
			l[i][j] = a[i][j]
		}
		for j in i .. n {
			u[i][j] = a[i][j]
		}
	}

	// Reconstruct PA = LU (apply permutation to original matrix)
	mut pa := original_a.clone()
	for i in 0 .. n {
		if ipiv[i] != i {
			// Swap rows i and ipiv[i]
			for j in 0 .. n {
				tmp := pa[i][j]
				pa[i][j] = pa[ipiv[i]][j]
				pa[ipiv[i]][j] = tmp
			}
		}
	}

	lu_product := matrix_multiply(l, u)
	assert nearly_equal_matrix(pa, lu_product, test_tolerance), 'getrf: PA != LU'
}

fn test_getri_basic() {
	// TODO: fix this test
	$if false {
		// Test matrix inversion
		mut a := [[4.0, 3.0], [3.0, 2.0]] // Well-conditioned 2x2
		original_a := a.clone()

		// Get LU factorization
		mut ipiv := getrf(mut a) or {
			assert false, 'getrf failed for getri test'
			return
		}

		// Compute inverse
		getri(mut a, mut ipiv) or { assert false, 'getri failed on 2x2 matrix' }

		// Check A * A^(-1) = I
		identity_check := matrix_multiply(original_a, a)
		expected_identity := create_identity(2)
		assert nearly_equal_matrix(identity_check, expected_identity, test_tolerance), 'getri: A * A^(-1) != I'

		// Check A^(-1) * A = I
		identity_check2 := matrix_multiply(a, original_a)
		assert nearly_equal_matrix(identity_check2, expected_identity, test_tolerance), 'getri: A^(-1) * A != I'
	}
}

// ============================================================================
// POTRF Tests - Cholesky Factorization
// ============================================================================

fn test_potrf_basic() {
	// Test 1: Simple 2x2 SPD matrix
	mut a := [[4.0, 2.0], [2.0, 3.0]] // SPD matrix
	original_a := a.clone()

	potrf(mut a, blas.Uplo.upper) or { assert false, 'potrf failed on 2x2 SPD matrix' }

	// Extract upper triangular Cholesky factor
	mut u := [][]f64{len: 2, init: []f64{len: 2, init: 0.0}}
	for i in 0 .. 2 {
		for j in i .. 2 {
			u[i][j] = a[i][j]
		}
	}

	// Check U'U = A
	ut := matrix_transpose(u)
	reconstructed := matrix_multiply(ut, u)
	assert nearly_equal_matrix(reconstructed, original_a, test_tolerance), "potrf: U'U != A"

	// Test 2: Larger SPD matrix
	spd_matrix := create_spd_matrix(5, 123)
	mut a_large := spd_matrix.clone()
	original_large := spd_matrix.clone()

	potrf(mut a_large, blas.Uplo.upper) or { assert false, 'potrf failed on 5x5 SPD matrix' }

	// Extract upper triangular part and verify
	mut u_large := [][]f64{len: 5, init: []f64{len: 5, init: 0.0}}
	for i in 0 .. 5 {
		for j in i .. 5 {
			u_large[i][j] = a_large[i][j]
		}
	}

	ut_large := matrix_transpose(u_large)
	reconstructed_large := matrix_multiply(ut_large, u_large)
	assert nearly_equal_matrix(reconstructed_large, original_large, test_tolerance), "potrf: U'U != A for 5x5 matrix"
}

// ============================================================================
// GEEV Tests - General Eigenvalue Problem
// ============================================================================

fn test_geev_basic() {
	// Test 1: Simple 2x2 symmetric matrix (real eigenvalues)
	a := [[3.0, 1.0], [1.0, 3.0]]

	wr, wi, vl, vr := geev(a, .left_ev_compute, .right_ev_compute) or {
		assert false, 'geev failed on 2x2 symmetric matrix'
		return
	}

	// Check eigenvalues are real (wi should be zero)
	assert float64.tolerance(wi[0], 0.0, test_tolerance), 'geev: expected real eigenvalue'
	assert float64.tolerance(wi[1], 0.0, test_tolerance), 'geev: expected real eigenvalue'

	// For symmetric matrix, eigenvalues should be 4 and 2
	mut eigenvals := [wr[0], wr[1]]
	eigenvals.sort()
	assert float64.tolerance(eigenvals[0], 2.0, test_tolerance), 'geev: incorrect eigenvalue'
	assert float64.tolerance(eigenvals[1], 4.0, test_tolerance), 'geev: incorrect eigenvalue'

	// Test 2: Verify eigenvalue equation A*v = λ*v for right eigenvectors
	for i in 0 .. 2 {
		if float64.tolerance(wi[i], 0.0, test_tolerance) {
			// Real eigenvalue
			mut v := [vr[0][i], vr[1][i]]
			mut av := [0.0, 0.0]

			// Compute A*v
			for j in 0 .. 2 {
				for k in 0 .. 2 {
					av[j] += a[j][k] * v[k]
				}
			}

			// Compute λ*v
			mut lv := [wr[i] * v[0], wr[i] * v[1]]

			assert float64.tolerance(av[0], lv[0], test_tolerance), 'geev: A*v != λ*v for eigenvalue ${i}'
			assert float64.tolerance(av[1], lv[1], test_tolerance), 'geev: A*v != λ*v for eigenvalue ${i}'
		}
	}
}

// ============================================================================
// SYEV Tests - Symmetric Eigenvalue Problem
// ============================================================================

fn test_syev_basic() {
	// Test 1: Simple 2x2 symmetric matrix
	mut a := [[3.0, 1.0], [1.0, 3.0]]
	original_a := a.clone()

	eigenvals := syev(mut a, .ev_compute, blas.Uplo.upper) or {
		assert false, 'syev failed on 2x2 symmetric matrix'
		return
	}

	// Check eigenvalues (should be 2 and 4 for this matrix)
	assert eigenvals.len == 2, 'syev: wrong number of eigenvalues'
	assert float64.tolerance(eigenvals[0], 2.0, test_tolerance), 'syev: incorrect first eigenvalue'
	assert float64.tolerance(eigenvals[1], 4.0, test_tolerance), 'syev: incorrect second eigenvalue'

	// Check that eigenvectors are orthonormal
	assert check_orthogonal(a, true), 'syev: eigenvectors not orthonormal'

	// Test 2: Verify eigenvalue equation A*V = V*D
	mut d := [][]f64{len: 2, init: []f64{len: 2, init: 0.0}}
	d[0][0] = eigenvals[0]
	d[1][1] = eigenvals[1]

	av := matrix_multiply(original_a, a) // A * V (V is stored in a after syev)
	vd := matrix_multiply(a, d) // V * D

	assert nearly_equal_matrix(av, vd, test_tolerance), 'syev: A*V != V*D'
}

// ============================================================================
// GEQRF/ORGQR Tests - QR Factorization
// ============================================================================

fn test_geqrf_orgqr() {
	// TODO: fix this test

	$if false {

		// Test QR factorization on various matrix sizes
		test_cases := [
			[3, 3], // Square matrix
			[5, 3], // Tall matrix
			[3, 5], // Wide matrix
		]

		for case in test_cases {
			m := case[0]
			n := case[1]

			// Create test matrix
			a_original := create_random_matrix(m, n, 456 + m + n)
			mut a := a_original.clone()

			// Compute QR factorization
			tau := geqrf(mut a) or {
				assert false, 'geqrf failed for ${m}x${n} matrix'
				return
			}

			// Extract R (upper triangular part)
			mut r := [][]f64{len: m, init: []f64{len: n, init: 0.0}}
			for i in 0 .. m {
				for j in i .. n {
					if j < n {
						r[i][j] = a[i][j]
					}
				}
			}

			// Generate Q using orgqr
			orgqr(mut a, tau) or { assert false, 'orgqr failed for ${m}x${n} matrix' }

			// Check that Q has orthonormal columns
			if m >= n {
				// For tall matrices, Q should have orthonormal columns
				qt := matrix_transpose(a)
				qtq := matrix_multiply(qt, a)
				identity_n := create_identity(n)
				assert nearly_equal_matrix(qtq, identity_n, ortho_tolerance), 'QR: Q not orthonormal for ${m}x${n}'
			}

			// Check QR = A_original (Q*R should reconstruct original matrix)
			qr_product := matrix_multiply(a, r)
			assert nearly_equal_matrix(qr_product, a_original, test_tolerance), 'QR: Q*R != A for ${m}x${n}'
		}

	}
}

// ============================================================================
// GESVD Tests - Singular Value Decomposition
// ============================================================================

fn test_gesvd_basic() {
	// TODO: fix this test
	$if false {
		// Test 1: Simple 3x2 matrix
		a := [[1.0, 2.0], [3.0, 4.0], [5.0, 6.0]]

		s, u, vt := gesvd(a, .svd_all, .svd_all) or {
			assert false, 'gesvd failed on 3x2 matrix'
			return
		}

		// Check dimensions
		assert s.len == 2, 'gesvd: wrong number of singular values'
		assert u.len == 3 && u[0].len == 3, 'gesvd: wrong U dimensions'
		assert vt.len == 2 && vt[0].len == 2, 'gesvd: wrong V^T dimensions'

		// Check that singular values are non-negative and sorted
		for i in 0 .. s.len - 1 {
			assert s[i] >= s[i + 1], 'gesvd: singular values not sorted'
			assert s[i] >= 0, 'gesvd: negative singular value'
		}

		// Check orthogonality: U^T * U = I and V^T * V = I
		assert check_orthogonal(u, true), 'gesvd: U not orthogonal'
		assert check_orthogonal(vt, false), 'gesvd: V^T not orthogonal'

		// Test 2: Reconstruct original matrix: A = U * Σ * V^T
		mut sigma := [][]f64{len: 3, init: []f64{len: 2, init: 0.0}}
		for i in 0 .. s.len {
			sigma[i][i] = s[i]
		}

		us := matrix_multiply(u, sigma)
		reconstructed := matrix_multiply(us, vt)

		assert nearly_equal_matrix(reconstructed, a, test_tolerance), 'gesvd: U*Σ*V^T != A'
	}
}

// ============================================================================
// Integration Tests - Combined Operations
// ============================================================================

fn test_integration_linear_system_methods() {
	// Test that different methods give same result for solving Ax = b
	n := 4
	a_orig := create_random_matrix(n, n, 789)

	// Make matrix well-conditioned by adding to diagonal
	mut a := a_orig.clone()
	for i in 0 .. n {
		a[i][i] += 5.0
	}

	b_orig := create_random_matrix(n, 1, 987)

	// Method 1: Direct solve with gesv
	mut a1 := a.clone()
	mut b1 := b_orig.clone()
	gesv(mut a1, mut b1) or { assert false, 'integration: gesv failed' }

	// Method 2: LU factorization + manual back-substitution would be more complex
	// For now, just verify the solution by substitution
	mut residual := matrix_multiply(a, b1)
	for i in 0 .. n {
		residual[i][0] -= b_orig[i][0]
	}
	residual_norm := matrix_norm(residual, 'fro')
	assert residual_norm < test_tolerance, 'integration: solution residual too large'
}

fn test_cholesky_vs_lu() {
	// For SPD matrices, both Cholesky and LU should work
	n := 3
	spd := create_spd_matrix(n, 654)
	b := create_random_matrix(n, 1, 321)

	// Solve with general LU (gesv)
	mut a_lu := spd.clone()
	mut b_lu := b.clone()
	gesv(mut a_lu, mut b_lu) or { assert false, 'cholesky vs LU: gesv failed' }

	// For Cholesky method, we'd need potrs (solve after potrf)
	// which isn't exposed in the current bindings
	// So just verify the LU solution is correct
	mut residual := matrix_multiply(spd, b_lu)
	for i in 0 .. n {
		residual[i][0] -= b[i][0]
	}
	residual_norm := matrix_norm(residual, 'fro')
	assert residual_norm < test_tolerance, 'cholesky vs LU: LU solution incorrect'
}

// ============================================================================
// Main Test Functions - Entry Points
// ============================================================================

fn test_lapack_basic_functionality() {
	test_gesv_basic()
	test_gesv_square_systems()
	test_getrf_basic()
	test_getri_basic()
}

fn test_lapack_advanced_functionality() {
	test_potrf_basic()
	test_geev_basic()
	test_syev_basic()
	test_geqrf_orgqr()
	test_gesvd_basic()
}

fn test_lapack_integration() {
	test_integration_linear_system_methods()
	test_cholesky_vs_lu()
}
