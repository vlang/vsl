
module quaternion

const (
	q_epsilon = (1e-14)
)
