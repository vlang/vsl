module noise
import math { abs }
import rand

const single_perlin_3d = f32(0.6107391600293113)

const cube_perlin_3d = [
	[
		[0.5, 0.5050048266819215, 0.5100372569900443],
		[0.49999512395332424, 0.5049999013347033, 0.5100322820703714],
		[0.49996196659450715, 0.5049664048058112, 0.5099984445007454]
	],
	[
		[0.5049950745885698, 0.5099997041643857, 0.5150313576483349],
		[0.5049901985418941, 0.5099947788181406, 0.5150263827306247],
		[0.504957041183077, 0.5099612822959435, 0.5149925451745017]
	],
	[
		[0.5099611901790586, 0.5149650429230547, 0.5199953367381234],
		[0.5099563141323828, 0.5149601175835047, 0.5199903618339162],
		[0.5099231567735657, 0.5149266211073663, 0.5199565243706847]
	]
]



fn test_perlin3d() {
    rand.seed([u32(114764230), 293925637])

    // Test single point
		// println(noise.perlin3d(0.125, 0.125, 0.125))
    assert abs(noise.perlin3d(0.125, 0.125, 0.125) - single_perlin_3d) < 1.0e-6

    // Test 3x3x3 grid
    for i in 0..3 {
        for j in 0..3 {
            for k in 0..3 {
                ii := i * 0.01
                jj := j * 0.01
                kk := k * 0.01
                assert abs(noise.perlin3d(f32(ii), f32(jj), f32(kk)) - cube_perlin_3d[i][j][k]) < 1.0e-6
            }
        }
    }
}
