module utils

import dl

pub const (
	default_paths = []string{}
)
