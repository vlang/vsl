module vsl

import vsl.quaternion
import vsl.consts
