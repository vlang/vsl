module lapack64
