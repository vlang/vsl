// Copyright (c) 2019-2020 Ulises Jeremias Cornejo Fandos. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.
module specfunc

const (
	a = [
		0.08333333333333333,
		-2.777777777777778e-3,
		7.936507936507937e-4,
		-5.952380952380952e-4,
		8.417508417508418e-4,
		-1.917526917526918e-3,
		6.410256410256410e-3,
		-0.02955065359477124,
		0.1796443723688307,
		-1.39243221690590
	]
)
