module vsl

pub const (
	version = '0.1'
)
