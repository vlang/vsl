// Copyright (c) 2019 Ulises Jeremias Cornejo Fandos. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.

module vsl

pub const (
	cgs_speed_of_light = 2.99792458e10 /* cm / s */
	cgs_gravitational_constant = 6.673e-8 /* cm^3 / g s^2 */
	cgs_plancks_constant_h = 6.62606896e-27 /* g cm^2 / s */
	cgs_plancks_constant_hbar = 1.05457162825e-27 /* g cm^2 / s */
	cgs_astronomical_unit = 1.49597870691e13 /* cm */
	cgs_light_year = 9.46053620707e17 /* cm */
	cgs_parsec = 3.08567758135e18 /* cm */
	cgs_grav_accel = 9.80665e2 /* cm / s^2 */
	cgs_electron_volt = 1.602176487e-12 /* g cm^2 / s^2 */
	cgs_mass_electron = 9.10938188e-28 /* g */
	cgs_mass_muon = 1.88353109e-25 /* g */
	cgs_mass_proton = 1.67262158e-24 /* g */
	cgs_mass_neutron = 1.67492716e-24 /* g */
	cgs_rydberg = 2.17987196968e-11 /* g cm^2 / s^2 */
	cgs_boltzmann = 1.3806504e-16 /* g cm^2 / k s^2 */
	cgs_molar_gas = 8.314472e7 /* g cm^2 / k mol s^2 */
	cgs_standard_gas_volume = 2.2710981e4 /* cm^3 / mol */
	cgs_minute = 6e1 /* s */
	cgs_hour = 3.6e3 /* s */
	cgs_day = 8.64e4 /* s */
	cgs_week = 6.048e5 /* s */
	cgs_inch = 2.54e0 /* cm */
	cgs_foot = 3.048e1 /* cm */
	cgs_yard = 9.144e1 /* cm */
	cgs_mile = 1.609344e5 /* cm */
	cgs_nautical_mile = 1.852e5 /* cm */
	cgs_fathom = 1.8288e2 /* cm */
	cgs_mil = 2.54e-3 /* cm */
	cgs_point = 3.52777777778e-2 /* cm */
	cgs_texpoint = 3.51459803515e-2 /* cm */
	cgs_micron = 1e-4 /* cm */
	cgs_angstrom = 1e-8 /* cm */
	cgs_hectare = 1e8 /* cm^2 */
	cgs_acre = 4.04685642241e7 /* cm^2 */
	cgs_barn = 1e-24 /* cm^2 */
	cgs_liter = 1e3 /* cm^3 */
	cgs_us_gallon = 3.78541178402e3 /* cm^3 */
	cgs_quart = 9.46352946004e2 /* cm^3 */
	cgs_pint = 4.73176473002e2 /* cm^3 */
	cgs_cup = 2.36588236501e2 /* cm^3 */
	cgs_fluid_ounce = 2.95735295626e1 /* cm^3 */
	cgs_tablespoon = 1.47867647813e1 /* cm^3 */
	cgs_teaspoon = 4.92892159375e0 /* cm^3 */
	cgs_canadian_gallon = 4.54609e3 /* cm^3 */
	cgs_uk_gallon = 4.546092e3 /* cm^3 */
	cgs_miles_per_hour = 4.4704e1 /* cm / s */
	cgs_kilometers_per_hour = 2.77777777778e1 /* cm / s */
	cgs_knot = 5.14444444444e1 /* cm / s */
	cgs_pound_mass = 4.5359237e2 /* g */
	cgs_ounce_mass = 2.8349523125e1 /* g */
	cgs_ton = 9.0718474e5 /* g */
	cgs_metric_ton = 1e6 /* g */
	cgs_uk_ton = 1.0160469088e6 /* g */
	cgs_troy_ounce = 3.1103475e1 /* g */
	cgs_carat = 2e-1 /* g */
	cgs_unified_atomic_mass = 1.660538782e-24 /* g */
	cgs_gram_force = 9.80665e2 /* cm g / s^2 */
	cgs_pound_force = 4.44822161526e5 /* cm g / s^2 */
	cgs_kilopound_force = 4.44822161526e8 /* cm g / s^2 */
	cgs_poundal = 1.38255e4 /* cm g / s^2 */
	cgs_calorie = 4.1868e7 /* g cm^2 / s^2 */
	cgs_btu = 1.05505585262e10 /* g cm^2 / s^2 */
	cgs_therm = 1.05506e15 /* g cm^2 / s^2 */
	cgs_horsepower = 7.457e9 /* g cm^2 / s^3 */
	cgs_bar = 1e6 /* g / cm s^2 */
	cgs_std_atmosphere = 1.01325e6 /* g / cm s^2 */
	cgs_torr = 1.33322368421e3 /* g / cm s^2 */
	cgs_meter_of_mercury = 1.33322368421e6 /* g / cm s^2 */
	cgs_inch_of_mercury = 3.38638815789e4 /* g / cm s^2 */
	cgs_inch_of_water = 2.490889e3 /* g / cm s^2 */
	cgs_psi = 6.89475729317e4 /* g / cm s^2 */
	cgs_poise = 1e0 /* g / cm s */
	cgs_stokes = 1e0 /* cm^2 / s */
	cgs_stilb = 1e0 /* cd / cm^2 */
	cgs_lumen = 1e0 /* cd sr */
	cgs_lux = 1e-4 /* cd sr / cm^2 */
	cgs_phot = 1e0 /* cd sr / cm^2 */
	cgs_footcandle = 1.076e-3 /* cd sr / cm^2 */
	cgs_lambert = 1e0 /* cd sr / cm^2 */
	cgs_footlambert = 1.07639104e-3 /* cd sr / cm^2 */
	cgs_curie = 3.7e10 /* 1 / s */
	cgs_roentgen = 2.58e-7 /* a s / g */
	cgs_rad = 1e2 /* cm^2 / s^2 */
	cgs_solar_mass = 1.98892e33 /* g */
	cgs_bohr_radius = 5.291772083e-9 /* cm */
	cgs_newton = 1e5 /* cm g / s^2 */
	cgs_dyne = 1e0 /* cm g / s^2 */
	cgs_joule = 1e7 /* g cm^2 / s^2 */
	cgs_erg = 1e0 /* g cm^2 / s^2 */
	cgs_stefan_boltzmann_constant = 5.67040047374e-5 /* g / k^4 s^3 */
	cgs_thomson_cross_section = 6.65245893699e-25 /* cm^2 */
)
