module vcl

#flag -I@VMODROOT

#include <vcl.h>
