module plot

// Font handles data to customize fonts
pub struct Font {
pub mut:
	color  string = 'black'
	family string = 'monospace'
	size   f64    = 16.
}
