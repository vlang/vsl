module vcl
