// Copyright (c) 2019 Ulises Jeremias Cornejo Fandos. All rights reserved.
// Use of this source code is governed by an MIT license
// that can be found in the LICENSE file.

module vsl

const(
	num_fine_structure = (7.297352533e-3) /* 1 */
	num_avogadro = (6.02214199e23) /* 1 / mol */
	num_yotta = (1e24) /* 1 */
	num_zetta = (1e21) /* 1 */
	num_exa = (1e18) /* 1 */
	num_peta = (1e15) /* 1 */
	num_tera = (1e12) /* 1 */
	num_giga = (1e9) /* 1 */
	num_mega = (1e6) /* 1 */
	num_kilo = (1e3) /* 1 */
	num_milli = (1e-3) /* 1 */
	num_micro = (1e-6) /* 1 */
	num_cml_nano = (1e-9) /* 1 */
	num_pico = (1e-12) /* 1 */
	num_femto = (1e-15) /* 1 */
	num_atto = (1e-18) /* 1 */
	num_zepto = (1e-21) /* 1 */
	num_yocto = (1e-24) /* 1 */
)
