module dl

import dl

pub const default_paths = []string{}
