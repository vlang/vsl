module lapack

import math
import vsl.blas

// dgetrf computes the LU decomposition of an m×n matrix A using partial
// pivoting with row interchanges.
//
// The LU decomposition is a factorization of A into
//
//	A = P * L * U
//
// where P is a permutation matrix, L is a lower triangular with unit diagonal
// elements (lower trapezoidal if m > n), and U is upper triangular (upper
// trapezoidal if m < n).
//
// On entry, a contains the matrix A. On return, L and U are stored in place
// into a, and P is represented by ipiv.
//
// ipiv contains a sequence of row interchanges. It indicates that row i of the
// matrix was interchanged with ipiv[i]. ipiv must have length min(m,n), and
// Dgetrf will panic otherwise. ipiv is zero-indexed.
//
// Dgetrf returns whether the matrix A is nonsingular. The LU decomposition will
// be computed regardless of the singularity of A, but the result should not be
// used to solve a system of equation.
pub fn dgetrf(m int, n int, mut a []f64, lda int, ipiv []int) {
	mn := math.min(m, n)

	if m < 0 {
		panic(m_lt0)
	}
	if n < 0 {
		panic(n_lt0)
	}
	if lda < math.max(1, n) {
		panic(bad_lda)
	}

	// quick return if possible
	if mn == 0 {
		return
	}

	if a.len < (m - 1) * lda + n {
		panic(short_a)
	}
	if ipiv.len < mn {
		panic(bad_len_ipiv)
	}

	nb := ilaenv(1, 'DGETRF', ' ', m, n, -1, -1)

	if nb <= 1 || nb >= mn {
		// use the unblocked algorithm.
		return dgetf2(m, n, mut a, lda, ipiv)
	}

	for j := 0; j < mn; j += nb {
		jb := math.min(mn - j, nb)

		// factor diagonal and subdiagonal blocks and test for exact singularity.
		dgetf2(m - j, jb, mut a[j * lda + j..], lda, ipiv[j..j + jb])

		for i := j; i <= math.min(m - 1, j + jb - 1); i++ {
			ipiv[i] += j
		}

		// apply interchanges to columns 1..j-1.
		dlaswp(j, mut a, lda, j, j + jb - 1, ipiv[..j + jb], 1)

		if j + jb < n {
			// apply interchanges to columns 1..j-1.
			mut slice := unsafe { a[j + jb..] }
			dlaswp(j, mut slice, lda, j, j + jb, ipiv[..j + jb], 1)

			blas.dtstrf(.left, .lower, .notrans, .unit, jb, n - j - jb, 1, a[j * lda + j..],
				lda, a[j * lda + j + jb..], lda)

			if j + jb < m {
				blas.dgemm(.notrans, .notrans, m - j - jb, n - j - jb, jb, -1, a[(j + jb) * lda + j..],
					lda, a[j * lda + j + jb..], lda, 1, a[(j + jb) * lda + j + jb..],
					lda)
			}
		}
	}
}
