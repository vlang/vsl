module vcl

#flag linux -lOpenCL
#flag windows -lOpenCL
#flag darwin -framework OpenCL
#flag -I@VMODROOT

#include <vcl.h>
