module vcldl

import dl

pub const (
	default_paths = []string{}
)
