module ml

fn test_init_forest() { assert 'init_forest' == 'init_forest'}
fn test_fit() { assert 'fit' == 'fit'}
fn test_predict() { assert 'predict' == 'predict'}