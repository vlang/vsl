module blas

#flag linux -O2 -I/usr/local/include -I/usr/lib -I@VROOT/blas
#flag linux -lopenblas -llapacke -L/usr/local/lib -L/usr/lib
#flag windows -O2
#flag windows -lopenblas -lgfortran
#flag darwin -I/usr/local/opt/openblas/include -I@VROOT/blas
#flag darwin -lopenblas -L/usr/local/opt/openblas/lib
