module consts
