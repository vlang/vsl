module vlas

#flag linux -O2 -I/usr/local/include -I/usr/lib
#flag linux -llapacke -L/usr/local/lib -L/usr/lib
#flag windows -O2
#flag windows -lopenblas -lgfortran
#flag darwin -I/usr/local/opt/openblas/include -I/usr/local/include
#flag darwin -llapacke -lopenblas -L/usr/local/opt/openblas/lib -L/usr/local/lib
#flag -I@VMODROOT
