module vcl

#flag linux -I@VMODROOT
#flag windows -I@VMODROOT
#flag darwin -I@VMODROOT

#include <vcl.h>
