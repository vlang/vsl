module vlas

#flag linux -O2 -I/usr/local/include -I/usr/lib
#flag linux -lopenblas -llapacke -L/usr/local/lib -L/usr/lib
#flag windows -O2
#flag windows -lopenblas -lgfortran
#flag darwin -I/usr/local/opt/openblas/include
#flag darwin -llapacke -lopenblas -L/usr/local/opt/openblas/lib
#flag -I@VMODROOT
